`default_nettype none

//  ┌─┐ ┌─┐ ┌─┐ ┌─┐ ┌─┐ ┌─┐ ┌─┐ ┌─┐ ┌─┐ ┌─┐ ┌─┐ ┌─┐ ┌─┐ ┌─┐ ┌─┐ ┌─┐ ┌─┐
// ─┘ └─┘ └─┘ └─┘ └─┘ └─┘ └─┘ └─┘ └─┘ └─┘ └─┘ └─┘ └─┘ └─┘ └─┘ └─┘ └─┘ └─ clk
//      ┌───────┐                   ┌───────────────────────┐
// ─────┘       └───────────────────┘                       └─────────── in
//          ┌───────┐                   ┌───────────────────────┐
// ─────────┘       └───────────────────┘                       └─────── past
//      ┌───┐                       ┌───┐
// ─────┘   └───────────────────────┘   └─────────────────────────────── rise
//              ┌───┐                                       ┌───┐
// ─────────────┘   └───────────────────────────────────────┘   └─────── fall

module edgedetect(in, rise, clk);

input in, clk;
output rise;

reg past;

always @(posedge clk) past <= in;

assign rise = in & !past;
//assign fall = !in & past;

endmodule

